module hazard_detector(
	input clock, reset,
	input [] 
	output [15:0] fowarding_data
	output to_foward_or_not);
	
	
	
	
endmodule

