module EXMEM_regi (
	input clock, 
	input reset, 
	input sw1_in, sw4_in, sw5_in,
	output reg sw1_out, sw4_out, sw5_out);
	
	always @(posedge clock or negedge reset) begin
		if (reset == 1'b0) begin
			sw1_out <= 1'b0;
			sw4_out <= 1'b0;
			sw5_out <= 1'b0;
		end else if (clock == 1'b1) begin
			sw1_out <= sw1_in;
			sw4_out <= sw4_in;
			sw5_out <= sw5_in;
		end
	end
	
endmodule
