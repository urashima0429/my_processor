module sixteen_to_twelve(
	input [15:0] in,
	output [11:0] out);

	assign out = in[11:0];
	
endmodule
